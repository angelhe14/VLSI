library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mivga is
	generic( constant h_pulse: integer := 96;
				constant h_bp: integer := 48;
				constant h_pixels: integer := 640;
				constant h_fp: integer := 16;
				constant v_pulse: integer := 2;
				constant v_bp: integer := 33;
				constant v_pixels: integer := 480;
				constant v_fp: integer := 10
	);
port( clk50Mhz: in std_logic;
		red: out std_logic_vector(3 downto 0);
		green: out std_logic_vector(3 downto 0);
		blue: out std_logic_vector(3 downto 0);
		h_sync: out std_logic;
		v_sync: out std_logic;
		dipsw: in std_logic_vector(3 downto 0);
		a,b,c,d,e,f,g: out std_logic);
end entity mivga;

architecture behavioral of mivga is
constant cero:   std_logic_vector(6 downto 0):= "0111111";
constant uno:    std_logic_vector(6 downto 0):= "0000110";
constant dos:    std_logic_vector(6 downto 0):= "1011011";
constant tres:   std_logic_vector(6 downto 0):= "1001111";
constant cuatro: std_logic_vector(6 downto 0):= "1100110";
constant cinco:  std_logic_vector(6 downto 0):= "1101101";
constant seis:   std_logic_vector(6 downto 0):= "1111101";
constant siete:  std_logic_vector(6 downto 0):= "0000111";
constant ocho:   std_logic_vector(6 downto 0):= "1111111";
constant nueve:  std_logic_vector(6 downto 0):= "1110011";
constant r1:   std_logic_vector(3 downto 0):= (OTHERS => '1');
constant r0:   std_logic_vector(3 downto 0):= (OTHERS => '0');
constant g1:   std_logic_vector(3 downto 0):= (OTHERS => '1');		
constant g0:   std_logic_vector(3 downto 0):= (OTHERS => '0');
constant b1:   std_logic_vector(3 downto 0):= (OTHERS => '1');
constant b0:   std_logic_vector(3 downto 0):= (OTHERS => '0');
--variable a,b,c,d,e,f: std_ logic;
signal conectornum: std_logic_vector(6 downto 0);
constant h_period: integer := h_pulse + h_bp + h_pixels + h_fp;
constant v_period: integer := v_pulse + v_bp + v_pixels + v_fp;
signal h_count: integer range 0 to h_period - 1 := 0;
signal v_count: integer range 0 to v_period - 1 := 0;
signal reloj_pixel: std_logic;
signal column: integer range 0 to h_period - 1 := 0;
signal row: integer range 0 to v_period - 1 := 0;
signal display_ena: std_logic;

begin

	relojpixel: process(clk50MHz) is
	begin
		if rising_edge(clk50MHz) then 
			reloj_pixel <= not reloj_pixel;
		end if;
	end process relojpixel;
	
	contadores: process(reloj_pixel)
	begin
		if rising_edge(reloj_pixel) then
			if h_count <(h_period-1) then
				h_count <= h_count + 1;
			else
				h_count <= 0;
				if v_count < (v_period - 1) then
					v_count <= v_count + 1;
				else
					v_count<= 0;
				end if;
			end if;
		end if;
	end process contadores;
	
	serial_hsync: process(reloj_pixel)
	begin
		if rising_edge(reloj_pixel) then 
			if h_count > (h_pixels + h_fp) or 
				h_count > (h_pixels + h_fp + h_pulse) then
				h_sync <= '0';
			else
				h_sync <= '1';
			end if;
		end if;
	end process serial_hsync;
	
	serial_vsync: process(reloj_pixel)
	begin
		if rising_edge(reloj_pixel) then 
			if v_count > (v_pixels + v_fp) or 
				v_count > (v_pixels + v_fp + v_pulse) then
				v_sync <= '0';
			else
				v_sync <= '1';
			end if;
		end if;
	end process serial_vsync;

	coords_pixel: process(reloj_pixel)
	begin
		if rising_edge(reloj_pixel) then
			if(h_count < h_pixels) then
				column <= h_count;
			end if;
			if(v_count < v_pixels) then
				row <= v_count;
			end if;
		end if;
	end process coords_pixel;

	display_enable: process(reloj_pixel)
	begin
		if rising_edge(reloj_pixel) then
			if(h_count < h_pixels and v_count < v_pixels) then
				display_ena <= '1';
			else
				display_ena <= '0';
			end if;
		end if;
	end process display_enable;
	
with (dipsw) select 
conectornum <=
					"0111111" when "0000",
					"0000110" when "0001",
					"1011011" when "0010",
					"1001111" when "0011",
					"1100110" when "0100",
					"1101101" when "0101",
					"1111101" when "0110",
					"0000111" when "0111",
					"1111111" when "1000",
					"1110011" when "1001",
					"0000000" when others;
	
	process (conectornum, row, column)
	begin
	case conectornum is
	when uno=>
		if((row>210 and row <240) and
		(column>140 and column<150)) then 
			red <= (others => '0');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>250 and row <280) and
		(column>140 and column<150)) then 
			red <= (others => '1');
			green <= (others => '0');
			blue <= (others => '0');
		else 
			red <= (others => '0');
			green <= (others => '0');
			blue <= (others => '0');
		end if;
			
	when dos=>
		if((row>200 and row <210) and
		(column>110 and column<140)) then 
			red <= (others => '0');
			green <= (others => '0');
			blue <= (others => '1');
		elsif((row>210 and row <240) and
		(column>140 and column<150)) then 
			red <= (others => '0');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>280 and row <290) and
		(column>110 and column<140)) then 
			red <= (others => '1');
			green <= (others => '1');
			blue <= (others => '1');
		elsif((row>250 and row <280) and
		(column>100 and column<110)) then 
			red <= (others => '0');
			green <= (others => '1');
			blue <= (others => '1');
		elsif((row>240 and row <250) and
		(column>110 and column<140)) then 
			red <= (others => '1');
			green <= (others => '0');
			blue <= (others => '1');	
		else 
			red <= (others => '0');
			green <= (others => '0');
			blue <= (others => '0');
		end if;
		
	when tres=>
		if((row>200 and row <210) and
		(column>110 and column<140)) then 
			red <= (others => '0');
			green <= (others => '0');
			blue <= (others => '1');
		elsif((row>210 and row <240) and
		(column>140 and column<150)) then 
			red <= (others => '0');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>250 and row <280) and
		(column>140 and column<150)) then 
			red <= (others => '1');
			green <= (others => '0');
			blue <= (others => '0');
		elsif((row>240 and row <250) and
		(column>110 and column<140)) then 
			red <= (others => '1');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>240 and row <250) and
		(column>110 and column<140)) then 
			red <= (others => '1');
			green <= (others => '0');
			blue <= (others => '1');	
		else 
			red <= (others => '0');
			green <= (others => '0');
			blue <= (others => '0');
		end if;

	when cuatro=>
		if((row>210 and row <240) and
		(column>140 and column<150)) then 
			red <= (others => '0');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>250 and row <280) and
		(column>140 and column<150)) then 
			red <= (others => '1');
			green <= (others => '0');
			blue <= (others => '0');
		elsif((row>210 and row <240) and
		(column>100 and column<110)) then 
			red <= (others => '1');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>240 and row <250) and
		(column>110 and column<140)) then 
			red <= (others => '1');
			green <= (others => '0');
			blue <= (others => '1');	
		else 
			red <= (others => '0');
			green <= (others => '0');
			blue <= (others => '0');
		end if;

	when cinco=>
		if((row>200 and row <210) and
		(column>110 and column<140)) then 
			red <= (others => '0');
			green <= (others => '0');
			blue <= (others => '1');
		elsif((row>280 and row <290) and
		(column>110 and column<140)) then 
			red <= (others => '0');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>250 and row <280) and
		(column>140 and column<150)) then 
			red <= (others => '1');
			green <= (others => '0');
			blue <= (others => '0');
		elsif((row>210 and row <240) and
		(column>100 and column<110)) then 
			red <= (others => '1');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>240 and row <250) and
		(column>110 and column<140)) then 
			red <= (others => '1');
			green <= (others => '0');
			blue <= (others => '1');	
		else 
			red <= (others => '0');
			green <= (others => '0');
			blue <= (others => '0');
		end if;

	when seis=>
		if((row>200 and row <210) and
		(column>110 and column<140)) then 
			red <= (others => '0');
			green <= (others => '0');
			blue <= (others => '1');
		elsif((row>250 and row <280) and
		(column>100 and column<110)) then 
			red <= (others => '0');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>280 and row <290) and
		(column>110 and column<140)) then 
			red <= (others => '0');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>250 and row <280) and
		(column>140 and column<150)) then 
			red <= (others => '1');
			green <= (others => '0');
			blue <= (others => '0');
		elsif((row>210 and row <240) and
		(column>100 and column<110)) then 
			red <= (others => '1');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>240 and row <250) and
		(column>110 and column<140)) then 
			red <= (others => '1');
			green <= (others => '0');
			blue <= (others => '1');	
		else 
			red <= (others => '0');
			green <= (others => '0');
			blue <= (others => '0');
		end if;
		
	when siete=>
		if((row>210 and row <240) and
		(column>140 and column<150)) then 
			red <= (others => '0');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>200 and row <210) and
		(column>110 and column<140)) then 
			red <= (others => '1');
			green <= (others => '0');
			blue <= (others => '0');
		elsif((row>250 and row <280) and
		(column>140 and column<150)) then 
			red <= (others => '1');
			green <= (others => '0');
			blue <= (others => '0');
		else 
			red <= (others => '0');
			green <= (others => '0');
			blue <= (others => '0');
		end if;
		
	when ocho=>
		if((row>200 and row <210) and
		(column>110 and column<140)) then 
			red <= (others => '0');
			green <= (others => '0');
			blue <= (others => '1');
		elsif((row>250 and row <280) and
		(column>100 and column<110)) then 
			red <= (others => '1');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>280 and row <290) and
		(column>110 and column<140)) then 
			red <= (others => '1');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>210 and row <240) and
		(column>140 and column<150)) then 
			red <= (others => '0');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>250 and row <280) and
		(column>140 and column<150)) then 
			red <= (others => '1');
			green <= (others => '0');
			blue <= (others => '0');
		elsif((row>210 and row <240) and
		(column>100 and column<110)) then 
			red <= (others => '1');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>240 and row <250) and
		(column>110 and column<140)) then 
			red <= (others => '1');
			green <= (others => '0');
			blue <= (others => '1');	
		else 
			red <= (others => '0');
			green <= (others => '0');
			blue <= (others => '0');
		end if;		

	when nueve=>
		if((row>200 and row <210) and
		(column>110 and column<140)) then 
			red <= (others => '0');
			green <= (others => '0');
			blue <= (others => '1');
		elsif((row>210 and row <240) and
		(column>140 and column<150)) then 
			red <= (others => '0');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>250 and row <280) and
		(column>140 and column<150)) then 
			red <= (others => '1');
			green <= (others => '0');
			blue <= (others => '0');
		elsif((row>210 and row <240) and
		(column>100 and column<110)) then 
			red <= (others => '1');
			green <= (others => '1');
			blue <= (others => '0');
		elsif((row>240 and row <250) and
		(column>110 and column<140)) then 
			red <= (others => '1');
			green <= (others => '0');
			blue <= (others => '1');	
		else 
			red <= (others => '0');
			green <= (others => '0');
			blue <= (others => '0');
		end if;
	end case;
	end process;
end architecture;